library verilog;
use verilog.vl_types.all;
entity send_control_vlg_vec_tst is
end send_control_vlg_vec_tst;
